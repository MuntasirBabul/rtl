`timescale 1ns/1ps

module tb_dual_port_ram();


