module axi_slave();

endmodule