`ifndef RAM_AGENT_PKG
`define RAM_AGENT_PKG

package ram_agent_pkg;
`include "uvm_macros.svh"
`include "ram_defines.svh"
`include "ram_seq_item.sv"
`include "ram_sequencer_0.sv"
`include "ram_sequencer_1.sv"
`include "ram_driver_0.sv"
`include "ram_driver_1.sv"
`include "ram_monitor_0.sv"
`include "ram_monitor_1.sv"
`include "ram_agent_0.sv"
`include "ram_agent_1.sv"
endpackage