class axi_common;
static mailbox gen2bfm = new();
endclass