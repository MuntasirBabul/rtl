class axi_mon;
task run();
    $display("#####_____ axi_mon _____#####");
endtask
endclass