class axi_cov;
task run();
    $display("#####_____ axi_cov _____#####");
endtask
endclass