`ifndef RAM_TEST_LIST
`define RAM_TEST_LIST

package ram_test_list;

import uvm_pkg::*
`include "uvm_macros.svh"

import ram_env_pkg::*
import ram_seq_list::*

`include "ram_test.sv"

endpackage
`endif