// interface components:
// ports, signals, modport and clocking block

interface axi_interface
(
    input logic clk,
    input logic rst
);
    


endinterface