// interface components:
// ports, signals, modport and clocking block

interface axi_interface();
    


endinterface